----------------------------------------------------------------------------------
-- Company:         Drone Infrastructure Inspection and Interaction (DIII) Group
-- Engineer:        Frederik Falk Nyboe
-- 
-- Create Date:     18/02/2022 13:51:00 AM
-- Design Name:     MagController
-- Module Name:     latch - Behavioral
-- Project Name:    PL-Mag-Sensor
-- Target Devices:  Ultra96-V2
-- Tool Versions:   2020.2
-- Description:    
-- 
-- Dependencies:    
-- 
-- Revision:
-- Revision         0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity latch is
    generic (
        n_bits  :   POSITIVE    :=  6
    );
    port(
        inp     :   in  STD_LOGIC_VECTOR(n_bits-1 downto 0);
		outp	:	out	STD_LOGIC_VECTOR(n_bits-1 downto 0) := (others => '0');
		q		:	in	STD_LOGIC
    );
end latch;

architecture Behavioral of latch is
begin
	process (q)
	begin
		if (q = '1') then
			outp <= inp;
		end if;
	end process;
end Behavioral;
